CDLv2�H�\                                		                                                        		      		                                                                                                                                                                      	           	                                                                                                                                                                                                                                                                                                                 	                                                	                                                                                                                                                                                                                 	                                                                                                                        	            	                                				                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            					       		         			                                      		                      	      	                                                                                                                                                                                                                                                                                                                                      				                                                                                                                                                                                                                                                  	                                      		                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 	                                                                                                                                                                                                                                                                                                                                                                                                                                                                 	                                                                    			                  	             				                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     	                               	                               		                                                                                                                                                                                                                                                                                                                                                  	                             	                                                                                                                                      	                                                                                                                                                  	                                                                          		  	                                                                                                                                                                                                                                                                                              	                                                                                                   	                                                                                                                                                       	                                                                                                                                                                                                                                                                                                                                                           	                                                                                                                                                                                                                                                                                                                                                                             	       	         	            			                   	                              		                         	                              	                                                            	                                                   					                                          	                                                                              	                                                                                                                                                                                                                                                    	           	                                                                                                                                   	                                                        	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  	                                                                                                                                            	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      	                                                                                                                           	                                                                                                     	            		                                                                           	                                                                                                                                                                                                                                                            			                                                                                                                                                                                                                                                                          		                   	 	                                                                                               	 		     	        	                                                                                                                                                                                                                       		                                                                           		                                                                                              		               	             		                                                                    				                                                                                                                                                                                                                                                                                                                                                                                                         		                                                                                                                                             	               	                                                                                                                                                                                                                                                                                                                                                                	                                                                                                                                                                                                                                                                                                                                                                                                                                              		          		                 	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     	                                                                                                                                   		                                	          	                  		                 					                    	  				       	         	        	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     